module not_gate(A, B);
	
	input A;
	output B;
	
	assign B = ~A;
	
endmodule